-- todo
-- data channel arbitrer
